-- |==== LIBRARIES =====|
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;		
USE STD.TEXTIO.ALL;					-- Entrada de datos por archivo
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_ArchivoDeRegistros IS
end TB_ArchivoDeRegistros;

ARCHITECTURE behaviour OF TB_ArchivoDeRegistros IS
	
	COMPONENT ArchivoDeRegistros
	PORT(
		--DATA_OUT : INOUT STD_LOGIC_VECTOR( 15 DOWNTO 0);
		SHAMT	: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		DIR	: IN STD_LOGIC;
		CLK	: IN STD_LOGIC;
		WR	: IN STD_LOGIC;
		
		-- MEMORIA RAM DISTRIBUIDA DE 3 PUERTOS
		ADDR_WR	: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		ADDR_RD1: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		ADDR_RD2: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		WD	: IN STD_LOGIC_VECTOR( 15 DOWNTO 0);
		DINOUT1	: INOUT STD_LOGIC_VECTOR( 15 DOWNTO 0);
		DOUT2	: OUT STD_LOGIC_VECTOR( 15 DOWNTO 0);
		SHE	: IN STD_LOGIC;  -- SHIFT ENABLE
		DIN	: INOUT STD_LOGIC_VECTOR( 15 DOWNTO 0);
	);
	END COMPONENT;
	
	
	--INPUTS
	SIGNAL SHAMT := STD_LOGIC_VECTOR( 3 DOWNTO 0) : = (OTHERS => '0');
	SIGNAL DIR := STD_LOGIC := '0';
	SIGNAL CLK := STD_LOGIC := '0';
	SIGNAL WR := STD_LOGIC := '0';
	
	SIGNAL ADDR_WR := STD_LOGIC_VECTOR( 3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL ADDR_RD1 := STD_LOGIC_VECTOR( 3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL ADDR_RD2 := STD_LOGIC_VECTOR( 3 DOWNTO 0) := (OTHERS => '0');
	
	SIGNAL WD := STD_LOGIC_VECTOR( 15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL SHE := STD_LOGIC := '0';
	
	--BiDirs
	SIGNAL DATA_OUT	: STD_LOGIC_VECTOR( 15 DOWNTO 0);
	SIGNAL DINOUT1 : STD_LOGIC_VECTOR( 15 DOWNTO 0);
	SIGNAL DIN : STD_LOGIC_VECTOR( 15 DOWNTO 0);
	
	--OUTPUTS
	SIGNAL DOUT2 : STD_LOGIC_VECTOR( 15 DOWNTO 0);
	
	--CLOCK : Se debe definir el tiempo por cada ciclo
	CONSTANT CLK_period : TIME := 10ns;
	
	
	
	
	
	
	
	
	
	
	
	