LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY BARREL_SHIFTER IS

	GENERIC(
		BUS_BARREL : INTEGER := 8
	);

	PORT(
		DATA_IN	: IN STD_LOGIC_VECTOR( BUS_BARREL - 1 DOWNTO 0);
		DATA_OUT: OUT STD_LOGIC_VECTOR( BUS_BARREL - 1 DOWNTO 0);
		SHIFT: IN STD_LOGIC_VECTOR( 2 DOWNTO 0);
		TYPE_SHIFT: IN STD_LOGIC		-- 1: Left Shifter , 0: Right Shifter
	); 
END BARREL_SHIFTER;

ARCHITECTURE BEHAVIOUR OF BARREL_SHIFTER IS
	BEGIN
		PSHIFT : PROCESS (SHIFT , DATA_IN)
		VARIABLE SHIFT_DATA : STD_LOGIC_VECTOR( BUS_BARREL - 1 DOWNTO 0);
		VARIABLE INDICE		: INTEGER RANGE -8 TO 7;
		
		BEGIN
			IF( TYPE_SHIFT = '1' ) THEN 	-- 1: Left Shifter
				SHIFT_DATA := DATA_IN;
				FOR	I IN 0 TO 2 LOOP
					FOR J IN 7 DOWNTO 0 LOOP
						IF( SHIFT(I) = '1' ) THEN
							INDICE := J - 2**I ;	
							IF( INDICE < 0 ) THEN	
								SHIFT_DATA( J ) := '0';
							ELSE
								SHIFT_DATA( J ) := SHIFT_DATA(INDICE);
							END IF;
						END IF;
					END LOOP;
				END LOOP;
				DATA_OUT <= SHIFT_DATA;
				
			ELSE						-- 0: Right Shifter
				SHIFT_DATA := DATA_IN;
				FOR	I IN 0 TO 2 LOOP
					FOR J IN 0 TO 7 LOOP
						IF( SHIFT(I) = '1' ) THEN
							INDICE := J + 2**I ;	
							IF( INDICE > 7 ) THEN	
								SHIFT_DATA( J ) := '0';
							ELSE
								SHIFT_DATA( J ) := SHIFT_DATA(INDICE);
							END IF;
						END IF;
					END LOOP;
				END LOOP;
				DATA_OUT <= SHIFT_DATA;
			END IF;
		END PROCESS PSHIFT;
	END BEHAVIOUR;

	