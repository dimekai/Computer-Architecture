library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity MEMORIA_PROGRAMA is
	PORT(
		A : in  STD_LOGIC_VECTOR (15 downto 0);
      D : out  STD_LOGIC_VECTOR (24 downto 0)
	);
end MEMORIA_PROGRAMA;

architecture MEMP of MEMORIA_PROGRAMA is
CONSTANT OPCODE_TIPOR 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000"; -- OPERACIONES _00 (TIPO R)
CONSTANT OPCODE_LI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
CONSTANT OPCODE_LWI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
CONSTANT OPCODE_SWI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
CONSTANT OPCODE_SW		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
CONSTANT OPCODE_ADDI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
CONSTANT OPCODE_SUBI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
CONSTANT OPCODE_ANDI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
CONSTANT OPCODE_ORI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
CONSTANT OPCODE_XORI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
CONSTANT OPCODE_NANDI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
CONSTANT OPCODE_NORI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
CONSTANT OPCODE_XNORI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
CONSTANT OPCODE_BEQI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
CONSTANT OPCODE_BNEI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
CONSTANT OPCODE_BLTI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
CONSTANT OPCODE_BLETI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";
CONSTANT OPCODE_BGTI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
CONSTANT OPCODE_BGETI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
CONSTANT OPCODE_B			: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";
CONSTANT OPCODE_CALL		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10100";
CONSTANT OPCODE_RET		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10101";
CONSTANT OPCODE_NOP		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10110";
CONSTANT OPCODE_LW 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10111";
--	FUNCONDE	
CONSTANT FUNCODE_ADD		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
CONSTANT FUNCODE_SUB		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
CONSTANT FUNCODE_AND		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
CONSTANT FUNCODE_OR		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
CONSTANT FUNCODE_XOR		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
CONSTANT FUNCODE_NAND	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
CONSTANT FUNCODE_NOR		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
CONSTANT FUNCODE_XNOR	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
CONSTANT FUNCODE_NOT		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
CONSTANT FUNCODE_SLL		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
CONSTANT FUNCODE_SRL		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
-- REGISTROS	
CONSTANT R0					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
CONSTANT R1					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
CONSTANT R2					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
CONSTANT R3					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
CONSTANT R4					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
CONSTANT R5					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
CONSTANT R6					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
CONSTANT R7					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
CONSTANT R8					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
CONSTANT R9					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
CONSTANT R10				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
CONSTANT R11				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1011";
CONSTANT R12				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100";
CONSTANT R13				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1101";
CONSTANT R14				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1110";
CONSTANT R15				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1111";
-- SIN USO	
CONSTANT SU					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";


TYPE ARR IS ARRAY (0 TO 2**16 - 1) OF STD_LOGIC_VECTOR(24 DOWNTO 0); 
CONSTANT ROM : ARR := (
		--CARGA DE NUMEROS
    opcode_LI & R0 & X"00E4", -- 10
    opcode_SWI & R0 & X"000A", -- 1
    opcode_LI & R0 & X"0032", -- 2
    opcode_SWI & R0 & X"000B", -- 3
    opcode_LI & R0 & X"FAD3", -- 8
    opcode_SWI & R0 & X"000C", -- 5
    opcode_LI & R0 & X"0204", -- 6
    opcode_SWI & R0 & X"000D", -- 7
    opcode_LI & R0 & X"F046", -- 4
    opcode_SWI & R0 & X"000E", -- 9
    opcode_LI & R0 & X"0017", -- 0
    opcode_SWI & R0 & X"000F", -- 11

	--i, j, limites
	opcode_LI & R0 & X"0000", -- 12
	opcode_LI & R1 & X"0000", -- 13
	opcode_LI & R2 & X"0000", -- 14
	opcode_LI & R3 & X"0006", -- 15

	--CICLO I
	opcode_SUBI & R4 & R3 & X"001", -- 16
	opcode_BGETI & R4 & R0 & X"00E", -- 17
	opcode_LI & R1 & X"0000", -- 18
	opcode_tipoR & R5 & R4 & R0 & SU & funcode_SUB, -- 19 
	opcode_BGETI & R5 & R1 & X"009", -- 20
	opcode_LW & R6 & R1 & X"00A", -- 21
	opcode_LW & R7 & R1 & X"00B", -- 22
	opcode_BLETI & R7 & R6 & X"004", -- 23
	opcode_LW & R2 & R1 & X"00A", -- 24
	opcode_SW & R7 & R1 & X"00A", -- 25
	opcode_SW & R2 & R1 & X"00B", -- 26
	opcode_ADDI & R1 & R1 & X"001", -- 27
	opcode_B & SU & X"0014", -- 28
	opcode_ADDI & R0 & R0 & X"001", -- 29
	opcode_B & SU & X"0011", -- 30
	opcode_NOP & SU & SU & SU & SU & SU, -- 31
	opcode_B & SU & X"001F", -- 32
		OTHERS=>(OTHERS=>'0')	--others para llenar de ceros las localidades y su tamaño.
);
begin
	D <= ROM( CONV_INTEGER(A) );
end MEMP;

