LIBRARY IEEE;
USE IEEE.library.STD_LOGIC_1164.ALL;
USE IEEE.library.STD_LOGIC_UNSIGNED.ALL;


--HACE CORRIMIENTO A LA DERECHA OPTIMIZADO

ENTITY BARRELS IS
	PORT (	DATAIN : in STD_LOGIC_VECTOR(7 DOWNTO 0);
			SHIFT  : in STD_LOGIC_VECTOR(2 DOWNTO 0);
			DATAOUT : out STD_LOGIC_VECTOR(7 DOWNTO 0)
		 );
end BARRELS;

ARCHITECTURE Behavioral OF BARRELS IS
	BEGIN
		PSSR : PROCESS ( DATAIN, SHIFT )
			DATAOUT <= TO_STDLOGICVECTOR(TO_BITVECTOR(DATAIN) SRL CONV_INTEGER(SHIFT));
	END PROCESS PSSR;
END Behavioral;
