-- |==== LIBRARIES =====|
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;		
USE STD.TEXTIO.ALL;					-- Entrada de datos
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_ArchivoDeRegistros IS
end TB_ArchivoDeRegistros;

ARCHITECTURE behaviour OF TB_ArchivoDeRegistros IS
	COMPONENT ArchivoDeRegistros
	PORT(
		--DATA_OUT : INOUT STD_LOGIC_VECTOR( 15 DOWNTO 0);
		SHAMT	: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		DIR		: IN STD_LOGIC;
		CLK 	: IN STD_LOGIC;
		WR		: IN STD_LOGIC;
		
		-- MEMORIA RAM DISTRIBUIDA DE 3 PUERTOS
		ADDR_WR	: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		ADDR_RD1: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		ADDR_RD2: IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
		WD		: IN STD_LOGIC_VECTOR( 15 DOWNTO 0);
		DINOUT1	: INOUT STD_LOGIC_VECTOR( 15 DOWNTO 0);
		DOUT2 	: OUT STD_LOGIC_VECTOR( 15 DOWNTO 0);
		SHE 	: IN STD_LOGIC;
				
	);