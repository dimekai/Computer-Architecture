LIBRARY IEEE;
USE IEEE.library.STD_LOGIC_1164.ALL;
USE IEEE.library.STD_LOGIC_UNSIGNED.ALL;


--HACE CORRIMIENTO A LA IZQUIERDA OPTIMIZADO

ENTITY BARRELS IS
	PORT (	DATAIN : in STD_LOGIC_VECTOR(7 DOWNTO 0);
			SHIFT  : in STD_LOGIC_VECTOR(2 DOWNTO 0);
			DATAOUT : out STD_LOGIC_VECTOR(7 DOWNTO 0)
		 );
end BARRELS;

ARCHITECTURE Behavioral OF BARRELS IS
	BEGIN
		PSSL : PROCESS ( DATAIN, SHIFT )
			DATAOUT <= TO_STDLOGICVECTOR(TO_BITVECTOR(DATAIN) SLL CONV_INTEGER(SHIFT));
	END PROCESS PSSL;
END Behavioral;
